//////////////////////////////////////////////////////////////////
//
// freqKeyMap.sv
// Anthony Nardomarino
// FPGA Piano Playing Robot
// MIT 6.111 Digital Systems Lab
// 11-15-2019
//
//////////////////////////////////////////////////////////////////

module freqKeyMap(
	input		[12:0]	freqIn,
	output	logic	[4:0]	keyOut
);
	logic	[4:0]	key;
	assign keyOut = key;
	always_comb begin
		case(freqIn)
			13'd7040: 	5'b11001;
			13'd6644: 	5'b11000;
			13'd6271: 	5'b10111;
			13'd5919: 	5'b10110;
			13'd5587: 	5'b10101;
			13'd5274: 	5'b10100;
			13'd4978: 	5'b10011;
			13'd4698: 	5'b10010;
			13'd4434: 	5'b10001;
			13'd4186: 	5'b10000;
			13'd3951: 	5'b11011;
			13'd3729: 	5'b11010;
			13'd3520: 	5'b11001;
			13'd3322: 	5'b11000;
			13'd3135: 	5'b10111;
			13'd2959: 	5'b10110;
			13'd2793: 	5'b10101;
			13'd2637: 	5'b10100;
			13'd2489: 	5'b10011;
			13'd2349: 	5'b10010;
			13'd2217: 	5'b10001;
			13'd2093: 	5'b10000;
			13'd1975: 	5'b11011;
			13'd1864: 	5'b11010;
			13'd1760: 	5'b11001;
			13'd1661: 	5'b11000;
			13'd1567: 	5'b10111;
			13'd1479: 	5'b10110;
			13'd1396: 	5'b10101;
			13'd1318: 	5'b10100;
			13'd1244: 	5'b10011;
			13'd1174: 	5'b10010;
			13'd1108: 	5'b10001;
			13'd1046: 	5'b10000;
			13'd987: 	5'b11011;
			13'd932: 	5'b11010;
			13'd880: 	5'b11001;
			13'd830: 	5'b11000;
			13'd783: 	5'b10111;
			13'd739: 	5'b10110;
			13'd698: 	5'b10101;
			13'd659: 	5'b10100;
			13'd622: 	5'b10011;
			13'd587: 	5'b10010;
			13'd554: 	5'b10001;
			13'd523: 	5'b10000;
			13'd493: 	5'b11011;
			13'd466: 	5'b11010;
			13'd440: 	5'b11001;
			13'd415: 	5'b11000;
			13'd391: 	5'b10111;
			13'd369: 	5'b10110;
			13'd349: 	5'b10101;
			13'd329: 	5'b10100;
			13'd311: 	5'b10011;
			13'd293: 	5'b10010;
			13'd277: 	5'b10001;
			13'd261: 	5'b10000;
			13'd246: 	5'b01011;
			13'd233: 	5'b01010;
			13'd220: 	5'b01001;
			13'd207: 	5'b01000;
			13'd195: 	5'b00111;
			13'd184: 	5'b00110;
			13'd174: 	5'b00101;
			13'd164: 	5'b00100;
			13'd155: 	5'b00011;
			13'd146: 	5'b00010;
			13'd138: 	5'b00001;
			13'd130: 	5'b00000;
			13'd123: 	5'b01011;
			13'd116: 	5'b01010;
			13'd110: 	5'b01001;
			13'd103: 	5'b01000;
			13'd97: 	5'b00111;
			13'd92: 	5'b00110;
			13'd87: 	5'b00101;
			13'd82: 	5'b00100;
			13'd77: 	5'b00011;
			13'd73: 	5'b00010;
			13'd69: 	5'b00001;
			13'd65: 	5'b00000;
			13'd61: 	5'b01011;
			13'd58: 	5'b01010;
			13'd55: 	5'b01001;
			13'd51: 	5'b01000;
			13'd48: 	5'b00111;
			13'd46: 	5'b00110;
		endcase
	end
endmodule // freqKeyMap

